library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bar_rom is
    port(
        clk: in std_logic;
        addr: in std_logic_vector(6 downto 0);
        data: out std_logic_vector(0 to 19)
    );
end bar_rom;

architecture content of bar_rom is
    type rom_type is array(0 to 127) of std_logic_vector(19 downto 0);
    constant BAR: rom_type :=
    (
        "11111101111111110111",
        "11010100000000010001",
        "10110010101010101101",
        "10011000100010000101",
        "10101000000000010011",
        "10101100000000000101",
        "10101100001000000101",
        "10100110001000000101",
        "10101110000101001011",
        "10100011010001010101",
        "10100101010000100101",
        "10100100101010100101",
        "10001001010100000101",
        "10100010001100000101",
        "10101000010110100011",
        "01001010010010010001",
        "10100000101110100111",
        "10100000000101010001",
        "10100000010010100111",
        "10100000000101100001",
        "10000010101011000111",
        "11100000001011000001",
        "10000010010110000111",
        "10100010001010000001",
        "10100001010100100111",
        "10100001010100100001",
        "10101010111000000111",
        "10100101101000010001",
        "10110111000000100111",
        "11011110000000100001",
        "10110000100001001011",
        "10101100000001000101",
        "10101000000100000101",
        "10101001000010000101",
        "10101000000000010101",
        "10100000000000000101",
        "10100000000000010011",
        "10100001000010010101",
        "10100000000001000101",
        "10100000000001000101",
        "11000000000100000011",
        "10100000000000000001",
        "10000010010000000111",
        "10100000010000000001",
        "10000000000000000111",
        "11100010001000000001",
        "10000100010000010111",
        "11100000000100000001",
        "10100010000000100111",
        "10110001000100010011",
        "10100010000001010101",
        "11011010000101000101",
        "10100000010100010011",
        "10010111010100010001",
        "10100001000001000111",
        "10100101110000000001",
        "10101010100000011111",
        "10101010110100000001",
        "11010001010000101011",
        "10101001011100000101",
        "10000100100000000101",
        "11100100101100000101",
        "10001001001000000101",
        "10100100100100010011",
        "10101000011000101011",
        "11010101001000101011",
        "10001000101010111011",
        "11100100101010001001",
        "10000001000000001011",
        "10100001010000001011",
        "10000000000000100111",
        "10100001000010010011",
        "10100100100001000111",
        "10100101000001010011",
        "10101000000000001111",
        "10100100000000001011",
        "10100000100000010111",
        "10100000100000101101",
        "10100000000001011011",
        "10100000000001010001",
        "10000000000010110111",
        "10101000000001100001",
        "10100000010110100101",
        "10100000001011000101",
        "10010000010111000011",
        "10101010011110000001",
        "10100010110000001111",
        "10100011110000000001",
        "10001001100000010111",
        "10100101100000010001",
        "10001011000000100111",
        "11001011000000000001",
        "10100110001000000111",
        "01010110000000000001",
        "10101000000001000111",
        "10101100000001000001",
        "10001100000000010111",
        "11101100000000000001",
        "10111000000000101011",
        "11011000000100000001",
        "10110000001000000111",
        "11111000000010000001",
        "10010000000100000101",
        "11011000010001000101",
        "10101000100010010011",
        "11011100000000000101",
        "10101100001000000101",
        "10100110001000000101",
        "10101110000101001011",
        "10100011010001010101",
        "10100101010000100101",
        "10100100101010100101",
        "10001001010100000101",
        "10100010001100000101",
        "10101000010110100011",
        "01001010010010010001",
        "10100000101110100111",
        "10100000000101010001",
        "10100000010010100111",
        "10100000000101100001",
        "10000010101011000111",
        "11100000001011000001",
        "10000010010110000111",
        "10100010001010000001",
        "10100001010100100111",
        "11010101011101010101",
        "10101101111010101111",
        "11111111111111111111"
    );
    signal addr_reg: std_logic_vector(6 downto 0);
begin
    process(clk)
    begin
        if clk'event and clk = '1' then
            addr_reg <= addr;
        end if;
    end process;            
    data <= BAR(conv_integer(addr_reg));
end content;

