library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity graphics is
end graphics;

architecture dispatcher of graphics is
begin

end dispatcher;