library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bar_rom is
    port(
        clk: in std_logic;
        addr: in std_logic_vector(5 downto 0);
        data: out std_logic_vector(0 to 19)
    );
end bar_rom;

architecture content of bar_rom is
    type rom_type is array(0 to 63) of std_logic_vector(19 downto 0);
    constant BAR: rom_type :=
    (
        "11111101111111110111",
        "11010100000000010001",
        "10110010101010101101",
        "10011000100010000101",
        "10101000000000010011",
        "10101100000000000101",
        "10101100001000000101",
        "10100110001000000101",
        "10101110000101001011",
        "10100011010001010101",
        "10100101010000100101",
        "10100100101010100101",
        "10001001010100000101",
        "10100010001100000101",
        "10101000010110100011",
        "01001010010010010001",
        "10100000101110100111",
        "10100000000101010001",
        "10100000010010100111",
        "10100000000101100001",
        "10000010101011000111",
        "11100000001011000001",
        "10000010010110000111",
        "10100010001010000001",
        "10100001010100100111",
        "10100001010100100001",
        "10101010111000000111",
        "10100101101000010001",
        "10110111000000100111",
        "11011110000000100001",
        "10110000100001001011",
        "10101100000001000101",
        "10001100000000010111",
        "11101100000000000001",
        "10111000000000101011",
        "11011000000100000001",
        "10110000001000000111",
        "11111000000010000001",
        "10010000000100000101",
        "11011000010001000101",
        "10101000100010010011",
        "11011100000000000101",
        "10101100001000000101",
        "10100110001000000101",
        "10101110000101001011",
        "10100011010001010101",
        "10100101010000100101",
        "10100100101010100101",
        "10001001010100000101",
        "10100010001100000101",
        "10101000010110100011",
        "01001010010010010001",
        "10100000101110100111",
        "10100000000101010001",
        "10100000010010100111",
        "10100000000101100001",
        "10000010101011000111",
        "11100000001011000001",
        "10000010010110000111",
        "10100010001010000001",
        "10100001010100100111",
        "11010101011101010101",
        "10101101111010101111",
        "11111111111111111111"
    );
    signal addr_reg: std_logic_vector(5 downto 0);
begin
    process(clk)
    begin
        if clk'event and clk = '1' then
            addr_reg <= addr;
        end if;
    end process;            
    data <= BAR(conv_integer(addr_reg));
end content;

